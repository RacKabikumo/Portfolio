`timescale 1ns/1ns
module Slt( in, out );
input in ;
output out ;

wire in, out ;


	assign out = in ;



endmodule