`timescale 1ns/1ns
module OR( dataA, dataB, out );
input dataA ;
input dataB ;
output out ;

wire dataA, dataB, out ;


	assign out = dataA | dataB ;



endmodule