`timescale 1ns/1ns
module AND( dataA, dataB, out );
input dataA ;
input dataB ;
output out ;

wire dataA, dataB, out ;

	and( out, dataA, dataB ) ;



endmodule